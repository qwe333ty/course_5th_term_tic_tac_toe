library ieee;
use ieee.std_logic_1164.all;

library work;
use work.game_utils.all;

entity MinMaxEngine is
end MinMaxEngine;

architecture MinMaxEngine_behaviour of MinMaxEngine is
    begin
end MinMaxEngine_behaviour;